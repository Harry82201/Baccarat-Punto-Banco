module tb_statemachine();

// Your testbench goes here. Make sure your tests exercise the entire design
// in the .sv file.  Note that in our tests the simulator will exit after
// 10,000 ticks (equivalent to "initial #10000 $finish();").

    logic slow_clock, resetb;
	logic [3:0] dscore, pscore, pcard3;
	logic load_pcard1, load_pcard2, load_pcard3;
    logic load_dcard1, load_dcard2, load_dcard3;
    logic player_win_light, dealer_win_light;
	
	statemachine STATEMACHINE (.*);
	
	initial begin
		slow_clock = 1'b0;
		forever #20 slow_clock = ~ slow_clock;
	end
	
	initial begin
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#10;
		assert(load_pcard1 == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		assert(load_dcard1 == 1);
		#80;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#10;
		assert(load_pcard2 == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#10;
		assert(load_dcard2 == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 7;
		#40;
		pscore = 8;
		#40;
		dscore = 5;
		#10;
		assert(load_pcard3 == 0);
		#40;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 8;
		#10;
		assert(load_pcard3 == 0);
		#40;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 9;
		#40;
		dscore = 8;
		#10;
		assert(load_pcard3 == 0);
		#40;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 9;
		#40;
		dscore = 9;
		#10;
		assert(load_pcard3 == 0);
		#40;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 6;
		#10;
		assert(load_pcard3 == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 7;
		#40;
		pcard3 = 8;
		pscore = 2;
		#10;
		assert(load_dcard3 == 0);
		#40;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 6;
		#40;
		pcard3 = 7;
		pscore = 1;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 5;
		#50;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 6;
		#40;
		pcard3 = 3;
		pscore = 7;
		#10;
		assert(load_dcard3 == 0);
		#40;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 5;
		#40;
		pcard3 = 7;
		pscore = 1;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 5;
		#50;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pcard3 = 3;
		pscore = 5;
		#10;
		assert(load_dcard3 == 0);
		#40;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 4;
		#40;
		pcard3 = 7;
		pscore = 1;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 1;
		#50;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 4;
		#40;
		pcard3 = 8;
		pscore = 2;
		#10;
		assert(load_dcard3 == 0);
		#40;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 3;
		#40;
		pcard3 = 7;
		pscore = 1;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 0;
		#50;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 3;
		#40;
		pcard3 = 8;
		pscore = 2;
		#10;
		assert(load_dcard3 == 0);
		#40;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 2;
		#40;
		pcard3 = 5;
		pscore = 9;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 5;
		#50;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 1;
		#40;
		pcard3 = 5;
		pscore = 9;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 9;
		#50;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 0;
		#40;
		pcard3 = 4;
		pscore = 8;
		#10;
		assert(load_dcard3 == 1);
		#30;
		dscore = 9;
		#50;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 7;
		#40;
		dscore = 2;
		#10;
		assert(load_pcard3 == 0);
		assert(load_dcard3 == 1);
		#30;
		dscore = 5;
		#50;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 7;
		#40;
		dscore = 2;
		#10;
		assert(load_pcard3 == 0);
		assert(load_dcard3 == 1);
		#30;
		dscore = 7;
		#50;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 7;
		#40;
		dscore = 2;
		#10;
		assert(load_pcard3 == 0);
		assert(load_dcard3 == 1);
		#30;
		dscore = 8;
		#50;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 7;
		#40;
		dscore = 6;
		#10;
		assert(load_pcard3 == 0);
		assert(load_dcard3 == 0);
		#40;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);
		#70;
		
		
		
		/*
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 3;
		#40;
		pscore = 7;
		#40;
		dscore = 9;
		#40;
		#10;
		assert(player_win_light == 0);
		assert(dealer_win_light == 1);//DWin
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 3;
		#40;
		pscore = 9;
		#40;
		dscore = 6;
		#40;
		#10;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);//PWin
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 3;
		#40;
		dscore = 6;
		#40;
		pscore = 9;
		#40;
		dscore = 8;
		#40; 
		#10;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);//PWin
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 1;
		#40;
		dscore = 0;
		#40;
		pscore = 9;
		#40;
		dscore = 9;
		#40; 
		#10;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);//Tie
		#70;
		
		resetb = 1'b0;
		#50;
		resetb = 1'b1;
		#40;
		pscore = 2;
		#40;
		dscore = 5;
		#40;
		pscore = 4;
		#40;
		dscore = 7;
		#40;
		pcard3 = 3;
		pscore = 7;
		#40;
		#10;
		assert(player_win_light == 1);
		assert(dealer_win_light == 1);//Tie
		#70;
		
		resetb = 1'b0;
		#40;
		resetb = 1'b1;
		#40;
		pscore = 4;
		#40;
		dscore = 5;
		#40;
		pscore = 1;
		#40;
		dscore = 6;
		#40;
		pcard3 = 8;
		pscore = 9;
		#40;
		#10;
		assert(player_win_light == 1);
		assert(dealer_win_light == 0);//Tie
		#70;
		*/
		
		$display("finished");
		
	end
						
endmodule

